// Code your testbench here
// or browse Examples
`include "driver.sv"
`include "intf.sv"
`include "tcm_mem_ram.v"
`include "tcm_mem.v"
`include "tb_top.v"