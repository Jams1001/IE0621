01101111
0
0
00100110
0
0
0
0
0
0
0
0
0
0
0
0