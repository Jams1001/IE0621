// Code your testbench here
// or browse Examples
`include "interface_1.sv"
`include "stimulus.sv"
`include "scoreboard.sv"
`include "reference_model.sv"
`include "driver.sv"
`include "monitor.sv"
`include "environment.sv"
`include "testcase.sv"
`include "tb_top.v"