`include "top_hvl.sv"
`include "interface.sv"
`include "reference_model.sv"
`include "driver.sv"
`include "monitor.sv"
`include "scoreboard.sv"
`include "agent.sv"
`include "env.sv"
`include "test_1.sv"
//`include "test_2.sv"
//`include "test_muldiv.sv"
`include "test_4.sv"
