// Code your testbench here
// or browse Examples
`include "stimulus.sv"
`include "interface_0.sv"
`include "interface_1.sv"
`include "driver.sv"
`include "monitor.sv"
`include "reference_model.sv"
`include "scoreboard.sv"
`include "environment.sv"
`include "testcase.sv"
`include "tb_top.v"
