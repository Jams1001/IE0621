// Code your design here
`include "uriscv_alu.v"
`include "uriscv_branch.v"
`include "uriscv_csr.v"
`include "uriscv_defs.v"
`include "uriscv_lsu.v"
`include "uriscv_muldiv.v"
`include "riscv_core.v"